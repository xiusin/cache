module cache

pub struct CacheOption {
}
